module my_and(
    input wire a, b,
    output wire c;
);
assign c = a & b
endmodule